--! @file spi_slave_tb.vhd
--!
--! @brief
--!
--! @copyright 2021 jstwinkles
--!
--! This program is free software: you can redistribute it and/or modify
--! it under the terms of the GNU General Public License as published by
--! the Free Software Foundation, either version 3 of the License, or
--! (at your option) any later version.
--!
--! This program is distributed in the hope that it will be useful,
--! but WITHOUT ANY WARRANTY; without even the implied warranty of
--! MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--! GNU General Public License for more details.
--!
--! You should have received a copy of the GNU General Public License
--! along with this program.  If not, see <https://www.gnu.org/licenses/>.

library ieee;
use ieee.std_logic_1164.all;

entity spi_slave_tb is
end spi_slave_tb;

architecture behavioral of spi_slave_tb is

  -----------
  -- Types --
  -----------

  ---------------
  -- Constants --
  ---------------

  -------------
  -- Signals --
  -------------

  -------------
  -- Aliases --
  -------------

begin

end behavioral;
